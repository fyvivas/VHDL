library verilog;
use verilog.vl_types.all;
entity codec_vlg_vec_tst is
end codec_vlg_vec_tst;
