library verilog;
use verilog.vl_types.all;
entity half_adder_vlg_vec_tst is
end half_adder_vlg_vec_tst;
